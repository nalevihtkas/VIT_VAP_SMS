module and(y,in2,in1);
input in1,in2;
output y;
assign y=in1&in2;
endmodule