module and_tb();

reg in1,in2;
wire y;

and ut(y,in2,in1);  

 initial 
 begin
 //test case 
 end
 endmodule